module mux_4 #(
    D_WIDTH = 32
)(
    input  logic [D_WIDTH-1:0] in0,
    input  logic [D_WIDTH-1:0] in1,
    input  logic [D_WIDTH-1:0] in2,
    input  logic [D_WIDTH-1:0] in3,
    input  logic [1:0]         sel,
    output logic [D_WIDTH-1:0] out
);
always_comb
case (sel)
    2'b00: out = in0;
    2'b01: out = in1;
    2'b10: out = in2;
    2'b11: out = in3;
    default: out = '0;
endcase

endmodule
