module pc_reg #(
    parameter WIDTH = 32
) (
    input  logic             clk,
    input  logic [WIDTH-1:0] pc_in,
    output logic [WIDTH-1:0] pc_out
);

always_ff @(posedge clk) begin
    pc_out <= pc_in;
end

endmodule
